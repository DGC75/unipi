module somma_differenza(output [N - 1: 0] out, output rip_out, input [N - 1: 0] inA, [N - 1: 0] inB);

    

endmodule