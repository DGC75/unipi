module testAdd2();
    


endmodule