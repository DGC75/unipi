//CONTATORE MOD4 DA 1bit
//PER OGNI VOLTA CHE VEDO UN 1, RESTITUIRE (cont++)%4
//IMPLEMENTAZIONE DI MEALY


module cntMod4(output [1:0]out, input in, input clk);
    


endmodule
    
