module s(output out, input inS, input in);
        xor(out, inS, in);
endmodule